module counter();
endmodule