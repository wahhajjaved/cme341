module basic_BCD_counter();
endmodule